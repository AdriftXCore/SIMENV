`ifndef __TOP_DEFINE_VH
`define __TOP_DEFINE_VH 1

`define DAT_W 32

`endif